module m1;
  logic [31:0] data;
  assign data = '0;
endmodule