module m1;
  logic [31:0] data;
  logic [31:0] data2;
  assign data = '0;
  assign data2 = '1;
endmodule